module vga_control_module
{
    
}